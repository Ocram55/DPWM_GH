`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:11:27 02/27/2016 
// Design Name: 
// Module Name:    Display 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Display(
	input wire [3:0] ones,tens,hundreds,mil,
	output wire [6:0] in0 ,in1,in2,in3
    );

reg [6:0] in00, in11,in22,in33;

// 7-segment encoding
//      0
//     ---
//  5 |   | 1
//     --- <--6
//  4 |   | 2
//     ---
//      3

   always @(ones)
      case (ones)
          4'b0001 : in00 = 7'b1111001;   // 1
          4'b0010 : in00 = 7'b0100100;   // 2
          4'b0011 : in00 = 7'b0110000;   // 3
          4'b0100 : in00 = 7'b0011001;   // 4
          4'b0101 : in00 = 7'b0010010;   // 5
          4'b0110 : in00 = 7'b0000010;   // 6
          4'b0111 : in00 = 7'b1111000;   // 7
          4'b1000 : in00 = 7'b0000000;   // 8
          4'b1001 : in00 = 7'b0010000;   // 9
          4'b1010 : in00 = 7'b0001000;   // A
          4'b1011 : in00 = 7'b0000011;   // b
          4'b1100 : in00 = 7'b1000110;   // C
          4'b1101 : in00 = 7'b0100001;   // d
          4'b1110 : in00 = 7'b0000110;   // E
          4'b1111 : in00 = 7'b0001110;   // F
          default : in00 = 7'b1000000;   // 0
      endcase

   always @(tens)
      case (tens)
          4'b0001 : in11 = 7'b1111001;   // 1
          4'b0010 : in11 = 7'b0100100;   // 2
          4'b0011 : in11 = 7'b0110000;   // 3
          4'b0100 : in11 = 7'b0011001;   // 4
          4'b0101 : in11 = 7'b0010010;   // 5
          4'b0110 : in11 = 7'b0000010;   // 6
          4'b0111 : in11 = 7'b1111000;   // 7
          4'b1000 : in11 = 7'b0000000;   // 8
          4'b1001 : in11 = 7'b0010000;   // 9
          4'b1010 : in11 = 7'b0001000;   // A
          4'b1011 : in11 = 7'b0000011;   // b
          4'b1100 : in11 = 7'b1000110;   // C
          4'b1101 : in11 = 7'b0100001;   // d
          4'b1110 : in11 = 7'b0000110;   // E
          4'b1111 : in11 = 7'b0001110;   // F
          default : in11 = 7'b1000000;   // 0
      endcase

   always @(hundreds)
      case (hundreds)
          4'b0001 : in22 = 7'b1111001;   // 1
          4'b0010 : in22 = 7'b0100100;   // 2
          4'b0011 : in22 = 7'b0110000;   // 3
          4'b0100 : in22 = 7'b0011001;   // 4
          4'b0101 : in22 = 7'b0010010;   // 5
          4'b0110 : in22 = 7'b0000010;   // 6
          4'b0111 : in22 = 7'b1111000;   // 7
          4'b1000 : in22 = 7'b0000000;   // 8
          4'b1001 : in22 = 7'b0010000;   // 9
          4'b1010 : in22 = 7'b0001000;   // A
          4'b1011 : in22 = 7'b0000011;   // b
          4'b1100 : in22 = 7'b1000110;   // C
          4'b1101 : in22 = 7'b0100001;   // d
          4'b1110 : in22 = 7'b0000110;   // E
          4'b1111 : in22 = 7'b0001110;   // F
          default : in22 = 7'b1000000;   // 0
      endcase
		
   always @(mil)
      case (mil)
          4'b0001 : in33 = 7'b1111001;   // 1
          4'b0010 : in33 = 7'b0100100;   // 2
          4'b0011 : in33 = 7'b0110000;   // 3
          4'b0100 : in33 = 7'b0011001;   // 4
          4'b0101 : in33 = 7'b0010010;   // 5
          4'b0110 : in33 = 7'b0000010;   // 6
          4'b0111 : in33 = 7'b1111000;   // 7
          4'b1000 : in33 = 7'b0000000;   // 8
          4'b1001 : in33 = 7'b0010000;   // 9
          4'b1010 : in33 = 7'b0001000;   // A
          4'b1011 : in33 = 7'b0000011;   // b
          4'b1100 : in33 = 7'b1000110;   // C
          4'b1101 : in33 = 7'b0100001;   // d
          4'b1110 : in33 = 7'b0000110;   // E
          4'b1111 : in33 = 7'b0001110;   // F
          default : in33 = 7'b1000000;   // 0
      endcase
		
assign in0=in00;
assign in1=in11;
assign in2=in22;
assign in3=in33;

endmodule
